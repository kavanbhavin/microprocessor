module adder(); // add all inputs and outputs inside parentheses

  // inputs
  
  
  // outputs
  
  
  // reg and internal variable definitions
  
  
  // implement module here

  
endmodule