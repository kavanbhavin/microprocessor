module shifter(A, LA, LR, Y, C); // add all inputs and outputs inside parentheses

  // inputs
  input [7:0] A;
  input LA;
  input LR;
  
  // outputs
  output [7:0] Y;
  output C;
  
  // reg and internal variable definitions
  
  
  // implement module here

  
endmodule