module cpu(CLK, RESET, EN_L, Iin, Din, PC, NextPC, DataA, DataB, DataC, DataD, MW);
  input         CLK;
  input         RESET;
  input         EN_L;
  input  [15:0] Iin;
  input  [7:0]  Din;
  
  output [7:0]  PC;
  output [7:0]  NextPC;
  output [7:0]  DataA;
  output [7:0]  DataB;
  output [7:0]  DataC;
  output [7:0]  DataD;
  output        MW;
  
  // comment the two lines out below if you use a submodule to generate PC/NextPC
  reg [7:0] PC;
  reg [7:0] NextPC;
  
  reg MW;
  
  
  
  // ADD YOUR CODE BELOW THIS LINE
  always @ (posedge CLK) begin
		if(RESET) PC <= 8'd0;
		else PC <= NextPC;
  end
  
  always@(*) begin
		//set NextPC to stuff here.
		
  end
  
  
  
  
  
  // ADD YOUR CODE ABOVE THIS LINE

endmodule